//`timescale 1ns / 1ps
`include "param.v"

module control_unit(
    input [31:0] instruction,
    input br_eq,
    input br_lt,
    output reg br_un,
    output reg npc_op,
    output reg rf_we,
    output reg [1:0]wb_sel,
    output reg [2:0] sext_op,
    output reg [3:0] alu_op,
    output reg [1:0]alua_sel,
    output reg [1:0]alub_sel,
    output reg dram_we,
    output reg rf_read_en   
    );
    wire [6:0] opcode;
    wire [2:0] fun3;
    wire [6:0] fun7;
    assign opcode=instruction[6:0];
    assign fun3=instruction[14:12];
    assign fun7=instruction[31:25];
    always @(*) begin
        case (opcode)
            `LW:begin
                br_un=0;
                npc_op=0;
                rf_we=1;
                wb_sel=2'b01;
                sext_op=`I;
                alu_op=`add;
                alua_sel=1;
                alub_sel=1;
                dram_we=0;
                rf_read_en=1;
            end
            `I_type:begin
                case (fun3)
                    `ADDI:begin
                        br_un=0;
                        npc_op=0;
                        rf_we=1;
                        wb_sel=2'b00;
                        sext_op=`I;
                        alu_op=`add;
                        alua_sel=1;
                        alub_sel=1;
                        dram_we=0;
                        rf_read_en=1;
                    end 
                    `SLLI:begin
                        br_un=0;
                        npc_op=0;
                        rf_we=1;
                        wb_sel=2'b00;
                        sext_op=`I;
                        alu_op=`sll;
                        alua_sel=1;
                        alub_sel=1;
                        dram_we=0;
                        rf_read_en=1;
                    end
                    `SLTI:begin
                        br_un=0;
                        npc_op=0;
                        rf_we=1;
                        wb_sel=2'b00;
                        sext_op=`I;
                        alu_op=`slt;
                        alua_sel=1;
                        alub_sel=1;
                        dram_we=0;
                        rf_read_en=1;
                    end
                    `SLTUI:begin
                        br_un=0;
                        npc_op=0;
                        rf_we=1;
                        wb_sel=2'b00;
                        sext_op=`I;
                        alu_op=`sltu;
                        alua_sel=1;
                        alub_sel=1;
                        dram_we=0;
                        rf_read_en=1;
                    end
                    `XORI:begin
                        br_un=0;
                        npc_op=0;
                        rf_we=1;
                        wb_sel=2'b00;
                        sext_op=`I;
                        alu_op=`logic_xor;
                        alua_sel=1;
                        alub_sel=1;
                        dram_we=0;
                        rf_read_en=1;
                    end
                    `I_rightshift:begin
                        if (fun7==`SRLI)begin
                            br_un=0;
                            npc_op=0;
                            rf_we=1;
                            wb_sel=2'b00;
                            sext_op=`I;
                            alu_op=`srl;
                            alua_sel=1;
                            alub_sel=1;
                            dram_we=0;
                            rf_read_en=1;
                        end
                        else if (fun7==`SRAI) begin
                            br_un=0;
                            npc_op=0;
                            rf_we=1;
                            wb_sel=2'b00;
                            sext_op=`I;
                            alu_op=`sra;
                            alua_sel=1;
                            alub_sel=1;
                            dram_we=0;
                            rf_read_en=1;
                        end                             
                    end
                    `ORI:begin
                        br_un=0;
                        npc_op=0;
                        rf_we=1;
                        wb_sel=2'b00;
                        sext_op=`I;
                        alu_op=`logic_or;
                        alua_sel=1;
                        alub_sel=1;
                        dram_we=0;
                        rf_read_en=1;
                    end
                    `ANDI:begin
                        br_un=0;
                        npc_op=0;
                        rf_we=1;
                        wb_sel=2'b00;
                        sext_op=`I;
                        alu_op=`logic_and;
                        alua_sel=1;
                        alub_sel=1;
                        dram_we=0;
                        rf_read_en=1;
                    end
                    default: begin 
                        br_un=0;
                        npc_op=0;
                        rf_we=0;
                        wb_sel=2'b00;
                        sext_op=`U;
                        alu_op=`add;               
                        alua_sel=0;
                        alub_sel=0;
                        dram_we=0;
                        rf_read_en=0;
                    end
                endcase
            end
            `SW:begin
                br_un=0;
                npc_op=0;
                rf_we=0;
                wb_sel=2'b00;
                sext_op=`S;
                alu_op=`add;
                alua_sel=1;
                alub_sel=1;
                dram_we=1;
                rf_read_en=1;
            end
            `R_type:begin
                case (fun3)
                    `R_algo:begin
                        if (fun7==`ADD)begin
                            br_un=0;
                            npc_op=0;
                            rf_we=1;
                            wb_sel=2'b00;
                            sext_op=`I;
                            alu_op=`add;
                            alua_sel=1;
                            alub_sel=0;
                            dram_we=0;
                            rf_read_en=1;
                        end
                        else if (fun7==`SUB) begin
                            br_un=0;
                            npc_op=0;
                            rf_we=1;
                            wb_sel=2'b00;
                            sext_op=`I;
                            alu_op=`sub;
                            alua_sel=1;
                            alub_sel=0;
                            dram_we=0;
                            rf_read_en=1;
                        end 
                    end 
                    `SLL:begin
                        br_un=0;
                        npc_op=0;
                        rf_we=1;
                        wb_sel=2'b00;
                        sext_op=`I;
                        alu_op=`sll;
                        alua_sel=1;
                        alub_sel=0;
                        dram_we=0;
                        rf_read_en=1;
                    end
                    `SLT:begin
                        br_un=0;
                        npc_op=0;
                        rf_we=1;
                        wb_sel=2'b00;
                        sext_op=`I;
                        alu_op=`slt;
                        alua_sel=1;
                        alub_sel=0;
                        dram_we=0;
                        rf_read_en=1;
                    end
                    `SLTU:begin
                        br_un=0;
                        npc_op=0;
                        rf_we=1;
                        wb_sel=2'b00;
                        sext_op=`I;
                        alu_op=`sltu;
                        alua_sel=1;
                        alub_sel=0;
                        dram_we=0;
                        rf_read_en=1;
                    end
                    
                    `XOR:begin
                        br_un=0;
                        npc_op=0;
                        rf_we=1;
                        wb_sel=2'b00;
                        sext_op=`I;
                        alu_op=`logic_xor;
                        alua_sel=1;
                        alub_sel=0;
                        dram_we=0;
                        rf_read_en=1;
                    end
                    `R_rightshift:begin
                        if (fun7==`SRL)begin
                            br_un=0;
                            npc_op=0;
                            rf_we=1;
                            wb_sel=2'b00;
                            sext_op=`I;
                            alu_op=`srl;
                            alua_sel=1;
                            alub_sel=0;
                            dram_we=0;
                            rf_read_en=1;
                        end
                        else if (fun7==`SRA) begin
                            br_un=0;
                            npc_op=0;
                            rf_we=1;
                            wb_sel=2'b00;
                            sext_op=`I;
                            alu_op=`sra;
                            alua_sel=1;
                            alub_sel=0;
                            dram_we=0;
                            rf_read_en=1;
                        end 
                    end
                    `OR:begin
                        br_un=0;
                        npc_op=0;
                        rf_we=1;
                        wb_sel=2'b00;
                        sext_op=`I;
                        alu_op=`logic_or;
                        alua_sel=1;
                        alub_sel=0;
                        dram_we=0;
                        rf_read_en=1;
                    end
                    `AND:begin
                        br_un=0;
                        npc_op=0;
                        rf_we=1;
                        wb_sel=2'b00;
                        sext_op=`I;
                        alu_op=`logic_and;
                        alua_sel=1;
                        alub_sel=0;
                        dram_we=0;
                        rf_read_en=1;
                    end
                    default: begin
                        br_un=0;
                        npc_op=0;
                        rf_we=0;
                        wb_sel=2'b00;
                        sext_op=`U;
                        alu_op=`add;               
                        alua_sel=0;
                        alub_sel=0;
                        dram_we=0;
                        rf_read_en=0;
                     end
                endcase
            end
            `LUI:begin
                br_un=0;
                npc_op=0;
                rf_we=1;
                wb_sel=2'b00;
                sext_op=`U;
                alu_op=`add;
                alua_sel=2;
                alub_sel=1;
                dram_we=0; 
                rf_read_en=0;
            end
            
            `AUIPC:begin
                br_un=0;
                npc_op=0;
                rf_we=1;
                wb_sel=2'b00;
                sext_op=`U;
                alu_op=`add;
                alua_sel=0;
                alub_sel=1;
                dram_we=0;
                rf_read_en=0;
            end
            `B_type:begin
                case (fun3)
                    `BEQ:begin
                        npc_op=br_eq;
                        rf_we=0;
                        wb_sel=2'b00;
                        sext_op=`B;
                        alu_op=`add;
                        alua_sel=0;
                        alub_sel=1;
                        dram_we=0;
                        br_un=0;
                        rf_read_en=1;
                    end 
                    `BNE:begin
                        npc_op=~br_eq;
                        rf_we=0;
                        wb_sel=2'b00;
                        sext_op=`B;
                        alu_op=`add;
                        alua_sel=0;
                        alub_sel=1;
                        dram_we=0;
                        br_un=0;
                        rf_read_en=1;
                    end
                    `BLT:begin
                        npc_op=br_lt;
                        rf_we=0;
                        wb_sel=2'b00;
                        sext_op=`B;
                        alu_op=`add;
                        alua_sel=0;
                        alub_sel=1;
                        dram_we=0;
                        br_un=0;
                        rf_read_en=1;
                    end
                    `BGE:begin
                        npc_op=~br_lt;
                        rf_we=0;
                        wb_sel=2'b00;
                        sext_op=`B;
                        alu_op=`add;
                        alua_sel=0;
                        alub_sel=1;
                        dram_we=0;
                        br_un=0;
                        rf_read_en=1;
                    end
                    `BLTU:begin
                        npc_op=br_lt;
                        rf_we=0;
                        wb_sel=2'b00;
                        sext_op=`B;
                        alu_op=`add;
                        alua_sel=0;
                        alub_sel=1;
                        dram_we=0;
                        br_un=1;
                        rf_read_en=1;
                    end
                    `BGEU:begin
                        npc_op=~br_lt;
                        rf_we=0;
                        wb_sel=2'b00;
                        sext_op=`B;
                        alu_op=`add;
                        alua_sel=0;
                        alub_sel=1;
                        dram_we=0;
                        br_un=1;
                        rf_read_en=1;
                    end
                    default: begin 
                        br_un=0;
                        npc_op=0;
                        rf_we=0;
                        wb_sel=2'b00;
                        sext_op=`U;
                        alu_op=`add;               
                        alua_sel=0;
                        alub_sel=0;
                        dram_we=0;
                        rf_read_en=0;
                    end
                endcase
            end
            `JARL:begin
                br_un=0;
                npc_op=1;
                rf_we=1;
                wb_sel=2'b10;
                sext_op=`I;
                alu_op=`add;
                alua_sel=1;
                alub_sel=1;
                dram_we=0;
                rf_read_en=1;
            end
            `JAL:begin
                br_un=0;
                npc_op=1;
                rf_we=1;
                wb_sel=2'b10;
                sext_op=`J;
                alu_op=`add;
                alua_sel=0;
                alub_sel=1;
                dram_we=0;
                rf_read_en=0;
            end
            default:begin 
                br_un=0;
                npc_op=0;
                rf_we=0;
                wb_sel=2'b00;
                sext_op=`U;
                alu_op=`add;               
                alua_sel=0;
                alub_sel=0;
                dram_we=0;
                rf_read_en=0;
            end 
        endcase
    end
endmodule
